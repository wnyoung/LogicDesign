
//���� ���� �ϴ� reset���� ��� �ϳ��� ���ľߵ�
module position_reset_n(	o_position_rst_n,
				i_sw0);

output	o_position_rst_n	;
input	i_sw0	;

assign o_position_rst_n = i_sw0;

endmodule